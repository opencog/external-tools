# vim:ts=20:
# swedish_phonet.dat - Swedish phonetic transformation rules for aspell
# Copyright (C) 2000  Martin Norb�ck  <d95mback@dtek.chalmers.se>
#
# This program is free software; you can redistribute it and/or
# modify it under the terms of the GNU General Public License
# as published by the Free Software Foundation; either version 2
# of the License, or (at your option) any later version.
# 
# This program is distributed in the hope that it will be useful,
# but WITHOUT ANY WARRANTY; without even the implied warranty of
# MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
# GNU General Public License for more details.
# 
# You should have received a copy of the GNU General Public License
# along with this program; if not, write to the Free Software
# Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA  02111-1307,
# USA.
#
# $Id: phonet.sv,v 1.2 2003/02/04 21:20:28 wobban Exp $
#
# ChangeLog:
# 2001-01-25: 0.2 total rewrite
# 2000-02-24: 0.1 initial version
#
# See end of file for description (in Swedish)

alphabet=[ABCDEFGHIJKLMNOPQRSTUVWXYZ���]

version 0.2

&	&
@	@
ANG(EIY��)-^	ANI	# f�rledet an- ska inte bli @-ljud
AGNO6	AKNO	# agnostiker osv.
AG(IE)-6	AK	# vokal+g(ie) ger ej j-ljud
A	A
BB-<	_
B	P
CCO-	K	# broccoli, piccolo
CC	KS	# successiv, access, succ�
CH	&	# choklad osv.
CK	K	# ck -> k som vanligt
C(EIY��)-<	S	# c + mjuk vokal -> s
C	K	# c + annat -> k
DJ(U��)-	I	# djungel, dj�vel, adj�
DD-	_
D	T
EG(IE)-6	EK	# vokal+g(ie) ger ej j-ljud
E	E
�	E
FF	F
F	F
G(EIY��)-3	I	# g+mjuk vokal ger j-ljud
GG6	K
GN	@N	# ugn, lugn...
G	K
H(AOU�EIY��)-^	H	# h i b�rjan av ord h�rs
H(AUO�EIY��)-	_	# annars stumt framf�r vokal
HJ	I	# hj->j (hj�rta osv.)
H	H
IG(IE)-6	IK	# vokal+g(ie) ger ej j-ljud
I	I
J	I
K(EIY��)-^	&	# k+mjuk vokal ger sje-ljud
KJ	&	# kjol
K	K
LJU-	I	# ljuga, ljus
LL-	_
L	L
MM-	_
M	M
NG6	@
NN-	_
N	N
ORIGI8	ORKI	# specialfall
OG(IE)-6	OK	# vokal+g(ie) ger ej j-ljud
O	O
PROJEKT	PRO&EKT	# specialfall
PSALT<	SALT	# specialfall
PSALM<	SALM	# specialfall
PP-	_
P	P
Q	K
RGI$6	RGI	# inget j i slutet
RGA$6	RIA	# h�r �r det d�remot j (arga,f�rga)
RGE$6	RIE	# h�r ocks� (Norge, �verge)
RGS$	RIS	# rgs i slutet
RG$	RI	# rg i slutet
RD	T	# "bl�tt" d
RN	N	# "bl�tt" n
RT	T	# "bl�tt" t
RLD	T	# v�rld
RL	L	# "bl�tt" l
RS	&	# sje-ljud (fars, g�rsg�rd)
RR-	_
R	R
SS-	_
SCHIZ6	SKITS	# specialfall
SCH6	&
SKJ	&	# skjorta, skjuta
SJ	&	# sje-ljud
S	S
TION9^	TION	# tionde
TION6	&ON	# station osv.
TT-	_
T	T
UG(IE)-6	UK	# vokal+g(ie) ger ej j-ljud
U	U
V	F
W	F
X9	KS
YG(IE)-6	YK	# vokal+g(ie) ger ej j-ljud
Y	I
ZZ	TS
Z	S
�TTIO9	OTIO	# specialfall (ej sje-ljud)
�RTION9	ORTION	# specialfall (r h�rs)
�G(IE)-6	OK	# vokal+g(ie) ger ej j-ljud
�	O
�G(IE)-6	EK	# vokal+g(ie) ger ej j-ljud
�	E
�G(IE)-6	�K	# vokal+g(ie) ger ej j-ljud
�	�

# Detta �r en lista med transformationer f�r att b�ttre kunna f�resl�
# ers�ttningsord till felstavade svenska ord.
#
# N�r man stavar fel p� grund av att man inte vet stavningen (till
# skillnad fr�n slarvfel), s� skriver man ofta n�got som skulle uttalas
# p� samma s�tt.
#
# F�r att kunna f�resl� b�ttre s� g�r aspell om ordet till en
# (ungef�rlig) fonetisk beskrivning med hj�lp av dessa regler.
#
# Det fungerar s� h�r:
#
# Ord som finns i ordlistan transformeras till sin fonetiska form
# N�r ett ord som inte finns med i ordlistan p�tr�ffas transformeras det
# till sin fonetiska form och j�mf�rs med de ord som finns i ordlistan.
# Det �r d�rf�r viktigt att ord som finns i ordlistan transformeras
# r�tt, annars kommer de aldrig att f�resl�s r�tt.
#
# F�ljande fonem finns:
# A kort och l�ngt a-ljud
# E kort och l�ngt e- och �-ljud
# F f- och v-ljud
# H tonande h (tonl�st h noteras inte)
# I kort och l�ngt i- och y-ljud, j-ljud
# K g- och k-ljud
# L l-ljud (�ven "bl�tt" som farlig och k�rl)
# M m-ljud
# N n-ljud (�ven "bl�tt" som barn och torn)
# O kort och l�ngt o- och �-ljud
# P b- och p-ljud
# R r-ljud
# S s-ljud
# T d- och t-ljud (�ven "bl�tt", som h�rd och h�rt)
# U u-ljud
# V v-ljud
# @ ng-ljud
# & sje-ljud
#
# S� h�r funkar transformeringsreglerna i korthet:
# * Det som st�r till v�nster transformeras till det till h�ger
# * St�r det ett eller flera - betyder det att de sista bokst�verna inte
#   �vers�tts, utan anv�nds n�sta g�ng
# * St�r det en siffra betyder det att den transformeringen har en viss
#   prioritet (normal prioritet �r 5), ju h�gre desto starkare
# * Inom varje initialbokstavsgrupp tilldelas prioritet uppifr�n och ner
#
# F�r mer information om processen och om aspell, se aspell.sourceforge.org
# Kapitel 5.3 i bruksanvisningen handlar om detta
